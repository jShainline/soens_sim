
B0 3 6 11 jjSFQ1 area=100
B1 3 8 12 jjSFQ1 area=100
B2 4 9 13 jjSFQ1 area=100
B3 5 10 14 jjSFQ1 area=100
 I0 0 2 pwl(0 0 1n 0 10n  22.78u )
 I1 0 3 pwl(0 0 0.09n 0 0.1n 265.00u )
I2 0 4 pwl(0 0 0.09n 0 0.1ns 0u)
 I3 0 5 pwl(0 0 0.09n 0 0.1ns  70.00u )
K1 L3 L4 1
 L0 3 4 20.60p 
L1 4 5 10.3p
L2 5 7 10.3n
L3 2 0 200p
L4 6 0 10.3p
L5 8 0 10.3p
L6 9 0 0.1f
L7 10 0 0.1f
R0 1 0 1
R1 7 0 R=v(1)+1e-6
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)
.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)

.control
set maxdata=2560000
tran 10p 102n
write ./dend_4jj_lin_ramp_100uA_Ide265.00uA_Isc070.00uA_Ljtl120.60pH.dat L2#branch v(5)
quit
.endc
